module top(
        input clk,
        input rst,
        input [31:0] inst
    );
    RegisterFile #(27, 32) rf

             endmodule
