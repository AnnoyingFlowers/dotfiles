module shift_rigister(

    );

endmodule
