module Decode #(INST_WIDTH = 1) (
        input [INST_WIDTH-1:0] inst,
        output imm,
        output rs1,
        output rs2,
        output rd
    );
endmodule
