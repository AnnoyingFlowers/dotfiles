module alu(

    );
endmodule
