module top(
        input clk,
        input rst,
        input [2:0] ctrl,
        input [8:0] in,
        output reg [8:0] out
    );

endmodule
