module shift_rigister(
        input clk,
        input rst,
        input in,
        output [7:0] out
    );

endmodule
