module alu(
        input [3:0] a,
        input [3:0] b,
        output [3:0] result,
        output carry,
        output zero,
        output overflow
    );
endmodule
