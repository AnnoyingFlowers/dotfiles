module shift_rigister(
        input clk,
        input rst,
        input in,
        output out,
        output [7:0] rigister
    );

endmodule
