module shift_rigister(
        input clk,
        input rst,
        input in,
        output out
    );

endmodule
