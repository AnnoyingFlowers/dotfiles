module key2ascii(
        input [7:0] key,
        output [7:0] ascii
    );
endmodule
