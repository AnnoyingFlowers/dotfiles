module shift_rigister(
        input clk,
        input rst,
        input [2:0] ctrl,
        input in,
        output [7:0] out
    );

    always @(posedge clk) begin
        ;
    end

endmodule
