module bcd7seg(
        input  [3:0] b,
        output reg [6:0] h
    );
    // detailed implementation ...

endmodule
