module alu(
        input [2:0] select,
        input [3:0] a,
        input [3:0] b,
        output [3:0] result,
        output carry,
        output zero,
        output overflow
    );
endmodule
