module barrel_shifter8(

    );
endmodule
