module top(
        input clk,
        input rst,
        input [31:0] inst,
        output reg [31:0] pc
    );
    wire [4:0] waddr;
    wire [31:0] wdata;
    wire wen;
    RegisterFile #(5, 32) R (
                     .clk(clk),
                     .waddr(waddr),
                     .wdata(wdata),
                     .wen(wen)
                 );
    Reg #(32, 32'x80000000)


    endmodule
