`timescale 1ns / 1ps
module kbd_ctrl(
        input clk,
        input rst,
        input ps2_clk,
        input ps2_data,
        output is_press,
        output [7:0] count,
        output [7:0] key
    );

    reg nextdata_n = 1'b1;
    reg [23:0] buffer;
    wire [7:0] count_reg = 8'b0;
    reg [7:0] current;
    wire [7:0] data;
    wire ready;
    wire overflow;

    ps2_keyboard u_ps2_keyboard(
                     .clk(clk),
                     .clrn(rst),
                     .ps2_clk(ps2_clk),
                     .ps2_data(ps2_data),
                     .nextdata_n(nextdata_n),
                     .data(data),
                     .ready(ready),
                     .overflow(overflow)
                 );

    key2ascii u_key2ascii(
                  .data   	( data ),
                  .ascii 	( current  )
              );

    always @(posedge clk) begin
        if(rst == 0) begin
            count_reg <= 8'b0;
            buffer <= 24'b0;
            nextdata_n <= 1'b1;
        end
        else begin
            if(nextdata_n == 1'b0)
                nextdata_n <= 1'b1;
            if(ready || overflow) begin
                if(current != 8'b0) begin
                    nextdata_n <= 1'b0;
                    buffer <= {buffer[15:0], current};
                end
            end
        end
    end

    assign is_press = (buffer[7:0] != 8'b0 && buffer[7:0] == buffer[15:8]) ? 1'b1 : 1'b0;

    always @(*) begin
        count_reg <= (buffer[15:8] == 8'hF0) ? count_reg + 1'b1 : count_reg;
    end

    assign count = count_reg;

    assign key = buffer[7:0];

endmodule
